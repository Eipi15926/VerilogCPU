module RF(wd,rr1,rr2,wr,rd1,rd2,clk,regwr);
    input[31:0] wd,rr1,rr2,wr,clk,regwr;
    output reg[31:0] rd1,rd2;

endmodule
//unused