module OR(oa,ob,oc);
input oa,ob;
output oc;
assign oc = oa|ob;
endmodule