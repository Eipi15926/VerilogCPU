module IM(addr,w,r,wd,rd);/*input : address in IM, output : instruction in address addr*/
    input [31:0] addr,wd;
    input w,r;
    output reg[31:0] rd;
    reg[31:0]Rom[31:0];//只是单纯地搬运了单周期的指令存储器IM并且没改名字，
    //并不是Read-Only Memory，是可读可写的正常存储器
    initial begin
        Rom[5'h00]=32'b000000_00001_00010_00000_00000_100000;//add $1,$2,$0
        Rom[5'h01]=32'b000000_00011_00010_00000_00000_100010;//sub
        Rom[5'h02]=32'b000000_00000_00001_00010_00000_100100;//and
        Rom[5'h03]=32'b000000_00000_00001_00010_00000_100101;//or
        Rom[5'h04]=32'b000000_00010_00011_00000_00000_101010;//slt
        //Rom[5'h05]=32'b000010_00000_00000_00000_00000_000000;//J 0
        Rom[5'h05]=32'b100011_00011_00000_0000_0000_0001_0000;//lw
        Rom[5'h06]=32'b101011_00011_00001_0000_0000_0001_0000;//sw
        Rom[5'h07]=32'b000100_00001_00010_1111_1111_1111_1110;//beq
        Rom[5'h08]=32'b000010_00000_00000_00000_00000_000000;//J 0
        //设以下为数据段
        Rom[5'h10]=32'h0321;
        Rom[5'h11]=32'h0;
    end
    always @(*)begin
        if (r)
            rd = Rom[addr[6:2]];
    end
    always @(*)begin
        if (w)
            Rom[addr[6:2]]=wd;
    end
endmodule
