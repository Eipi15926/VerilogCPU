module AND(br,aluz,mc);
input br,aluz;
output mc;
assign mc = br & aluz;
endmodule