module IM(addr,instr);/*input : address in IM, output : instruction in address addr*/
    input [31:0] addr;
    output [31:0] instr;
    wire[31:0]Rom[31:0];
        assign Rom[5'h00]=32'b000000_00001_00010_00000_00000_100000;//add $1,$2,$0
        assign Rom[5'h01]=32'b000000_00011_00010_00000_00000_100010;//sub
        assign Rom[5'h02]=32'b000000_00000_00001_00010_00000_100100;//and
        assign Rom[5'h03]=32'b000000_00000_00001_00010_00000_100101;//or
        assign Rom[5'h04]=32'b000000_00010_00011_00000_00000_101010;//slt
        //assign Rom[5'h05]=32'b000010_00000_00000_00000_00000_000000;//J 0
        assign Rom[5'h05]=32'b100011_00011_00000_0000_0000_0001_0000;//lw
        assign Rom[5'h06]=32'b101011_00011_00001_0000_0000_0001_0000;//sw
        assign Rom[5'h07]=32'b000100_00001_00010_1111_1111_1111_1110;//beq
        assign Rom[5'h08]=32'b000010_00000_00000_00000_00000_000000;//J 0
    assign instr = Rom[addr[6:2]];
endmodule
