module shl2(src,dst);
    input src[31:0];
    output dst[31:0];
endmodule